library verilog;
use verilog.vl_types.all;
entity ramSinglePort_vlg_vec_tst is
end ramSinglePort_vlg_vec_tst;
