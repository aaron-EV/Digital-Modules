library verilog;
use verilog.vl_types.all;
entity singlePort_ramSR_vlg_vec_tst is
end singlePort_ramSR_vlg_vec_tst;
