library verilog;
use verilog.vl_types.all;
entity modM_counter_vlg_vec_tst is
end modM_counter_vlg_vec_tst;
