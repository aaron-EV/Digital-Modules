library verilog;
use verilog.vl_types.all;
entity singlePort_ramRA_vlg_vec_tst is
end singlePort_ramRA_vlg_vec_tst;
