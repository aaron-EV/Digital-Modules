library verilog;
use verilog.vl_types.all;
entity \register\ is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        inReg           : in     vl_logic_vector(7 downto 0);
        outReg          : out    vl_logic_vector(7 downto 0)
    );
end \register\;
