library verilog;
use verilog.vl_types.all;
entity dualPort_ramSR_vlg_vec_tst is
end dualPort_ramSR_vlg_vec_tst;
