library verilog;
use verilog.vl_types.all;
entity modN_counter_vlg_vec_tst is
end modN_counter_vlg_vec_tst;
