library verilog;
use verilog.vl_types.all;
entity swapper_vlg_vec_tst is
end swapper_vlg_vec_tst;
